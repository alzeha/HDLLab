//Verilog HDL for "HDL_lab", "And" "functional"


module And (a, b, c);

	input a, b;
	output c;

	assign c = a && b;

endmodule
