//Verilog HDL for "HDL_lab", "one" "functional"


module one (out );

	output out;

	assign out = 1'b1;

endmodule
